/home/viterbi/09/lijunlia/work_gpdk045/LVS/netlist